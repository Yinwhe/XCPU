`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    21:34:44 03/12/2012
// Design Name:
// Module Name:    REGS ID/EX Latch
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module    REG_ID_EX(input clk,                                         //ID/EX Latch
                    input rst,
                    input EN,                                          //�?水�??�??�使�??
                    input flush,                                       //?��??�?�?�??�并�?�?�?DStall
                    input [31:0] IR_ID,                                //�???�?????�?(�?�?)
                    input [31:0] PCurrent_ID,                          //�???�?????令�???��?��??�??
                    input [4:0] rs1_addr,                               //�?????令�?��?��??�???A?��??
                    input [4:0] rs2_addr,                               //�?????令�?��?��??�???B?��??
                    input [31:0] rs1_data,                             //�?????令�?��?��??�???A?��??
                    input [31:0] rs2_data,                             //�?????令�?��?��??�???A?��??
                    input [31:0] Imm32,                                //�?????令�?��?�并?��?32�?�??��?��?
                    input [4:0]  rd_addr,                              //�?????令�?��?��??????�??��?��?
                    input ALUSrc_A,                             //�?????令�????�?ALU A?????��??
                    input ALUSrc_B,                             //�?????令�????�?ALU B?????��??
                    input [3:0]  ALUC,                                 //�?????令�????�?ALU??�??��??
                    input DatatoReg,                            //�?????令�????�?REG???��??�??��??????
                    input RegWrite,                                    //�?????令�????�?�?�??��??信�?
                    input WR,                                          //�?????令�????�?�??��?��?��??信�??
                    input [2:0] u_b_h_w,
                    input MIO,

                    output reg[31:0] PCurrent_EX,                      //??�?�???�?????令�?��??
                    output reg[31:0] IR_EX,                            //??�?�???�?????�?(�?�?)
                    output reg[4:0]  rs1_EX,
                    output reg[4:0]  rs2_EX,
                    output reg[31:0] A_EX,                             //??�?�???�?????令�?��?��??�???A?��??
                    output reg[31:0] B_EX,                             //??�?�???�?????令�?��?��??�???B?��??
                    output reg[31:0] Imm32_EX,                          //??�?�???�?????�?32�?�??��?��?
                    output reg[4:0]  rd_EX,                            //??�?�???�?????令�??????�?�??��?��??
                    output reg       ALUSrc_A_EX,                      //??�?�???�?????�?ALU A?????��??
                    output reg       ALUSrc_B_EX,                      //??�?�???�?????�?ALU B?????��??(�???)
                    output reg[3:0]  ALUC_EX,                          //??�?�???�?????�?ALU??�????��?��??
                    output reg       DatatoReg_EX,                     //??�?�???�?????�?REG???��??�??��??????
                    output reg       RegWrite_EX,                      //??�?�???�?????令�??�??��??信�??
                    output reg       WR_EX,                            //??�?�???�?????令�???��?��?��??信�?
                    output reg[2:0]  u_b_h_w_EX,
                    output reg       MIO_EX
                );

    always @(posedge clk or posedge rst) begin                           //ID/EX Latch
    if(rst) begin
        rd_EX        <= 0;
        RegWrite_EX  <= 0;
        WR_EX        <= 0;
        IR_EX        <= 32'h00000000;
        PCurrent_EX  <= 32'h00000000 ;
        rs1_EX       <= 0;
        rs2_EX       <= 0;
        MIO_EX       <= 0;
    end
    else if(EN)begin
            if(flush)begin                               //?��???��???��?��?��?水线�?止�?��??CPU?��??
                IR_EX       <= 32'h00000000;             //nop,�?�?�??????? : ????32'h00000013
                rd_EX       <= 0;                        //cancel Instruction write address
                RegWrite_EX <= 0;                        //�?�??��??信�?��?�?止�??�???�??
                WR_EX       <= 0;                        //cancel write memory
                PCurrent_EX <= PCurrent_ID;              //�?�??�?PC(�?�?)
                MIO_EX       <= 0;
            end
            else begin                                   //???��???��??正常�?�???EX�??
                PCurrent_EX <= PCurrent_ID;              //�?�??��?????令�?��?
                IR_EX       <= IR_ID;                    //�?�??��?????令�?��?(�?�?)
                A_EX        <= rs1_data;                 //�?�??��??�???A读�?��?��??
                B_EX        <= rs2_data;                 //�?�??��??�???B读�?��?��??
                Imm32_EX    <= Imm32;                    //�?�??��?��???�??��?
                rd_EX       <= rd_addr;                  //�?�??��??????�?�??��?��?
                rs1_EX      <= rs1_addr;
                rs2_EX      <= rs2_addr;
                ALUSrc_A_EX <= ALUSrc_A;                 //�?�??�?ALU A?????��?�信??
                ALUSrc_B_EX <= ALUSrc_B;                 //�?�??�?ALU B?????��?�信??
                ALUC_EX     <= ALUC;                     //�?�??�?ALU??�????��?��?�信??
                DatatoReg_EX<= DatatoReg;               //�?�??�?REG???��??�??��??????
                RegWrite_EX <= RegWrite;                 //�?�??��??�??��??信�?
                WR_EX       <= WR;                       //�?�??��???��?��?��??信�??
                u_b_h_w_EX    <= u_b_h_w;
                MIO_EX       <= MIO;

                end
        end
    end

endmodule